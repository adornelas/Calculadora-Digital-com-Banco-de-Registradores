module LetraE (
	output [6:0] Out
);

assign Out = ~7'b1111001;
endmodule