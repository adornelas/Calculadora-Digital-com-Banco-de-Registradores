module LetraO (
	output [6:0] Out
);

assign Out = ~7'b1011100;
endmodule