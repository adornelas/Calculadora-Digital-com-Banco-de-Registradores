module LetraR (
	output [6:0] Out
);

assign Out = ~7'b1010000;
endmodule